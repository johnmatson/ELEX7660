module seqDetect (  output logic valid,
                    input logic a, input logic [3:0] seq,
                    input logic clk, reset_n);

endmodule