module shiftReg #(parameter N = 8) (output logic [N-1:0] q,
                                    input logic [N-1:0] a,
                                    input logic [1:0] s
                                    input logic shiftIn, clk, reset_n);

endmodule