module vendingMachine ( output logic valid,
                        input logic nichel, dime, quarter,
                        input logic clk, reset_n);

endmodule