
module lab4 (
	clk_clk,
	led_export,
	reset_reset_n,
	spkr_export);	

	input		clk_clk;
	output	[7:0]	led_export;
	input		reset_reset_n;
	output		spkr_export;
endmodule
